LFSR/LFSR.sv