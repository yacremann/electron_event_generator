lookup_table_spectrum/LUT_spectrum.sv